* No part of this file can be released without the consent of SMIC.
* 
************************************************************************************  
*          NWell resistor under STI subcircuit netlist                             *  
************************************************************************************ 
.subckt rnwsti_ckt n2 n1 sub l=lr w=wr  
.param  
+rsh      = '653.4+drsh_rnwsti'   rtc1   = 8.36E-04       rtc2 = 9.42E-06   
+dw       = '1.28E-07+ddw_rnwsti'  
*+vc1     = 1.33E-02                vc2   = -4.64E-04  
+jc1a     = -1.80E-03              jc1b   = 2.66E-07    
+jc2a     = 8.27E-10               jc2b   = -9.83E-14
+rvc1     = 'jc1a+jc1b/l'          rvc2   = '(jc2a+jc2b/l)/l' 
+weff     = 'w-2*dw' 
+tcoef(temper)     = '1.0+(temper-25.0)*(rtc1+rtc2*(temper-25.0))' 

D1    sub  n2 nwdioll area='weff*l/5' pj='weff+2*l/5'
R1    n2   na 'rsh*l/4/weff*tcoef(temper)*min(max(1.0+rvc1*v(n2,n1)+rvc2*v(n2,n1)*v(n2,n1), 0.85), 1.15)' 
D2    sub  na nwdioll area='weff*l/5' pj='2*l/5'
R2    na   nb 'rsh*l/4/weff*tcoef(temper)*min(max(1.0+rvc1*v(n2,n1)+rvc2*v(n2,n1)*v(n2,n1), 0.85), 1.15)' 
D3    sub  nb nwdioll area='weff*l/5' pj='2*l/5'
R3    nb   nc 'rsh*l/4/weff*tcoef(temper)*min(max(1.0+rvc1*v(n2,n1)+rvc2*v(n2,n1)*v(n2,n1), 0.85), 1.15)' 
D4    sub  nc nwdioll area='weff*l/5' pj='2*l/5'
R4    nc   n1 'rsh*l/4/weff*tcoef(temper)*min(max(1.0+rvc1*v(n2,n1)+rvc2*v(n2,n1)*v(n2,n1), 0.85), 1.15)' 
D5    sub  n1 nwdioll area='weff*l/5' pj='weff+2*l/5'  
.ends rnwsti_ckt  
************************************************************************************  
*           NWell resistor under AA subcircuit netlist                             *  
************************************************************************************ 
.subckt rnwaa_ckt n2 n1 sub l=lr w=wr  
.param  
+rsh      = '373.00+drsh_rnwaa'    rtc1   = 1.77E-03       rtc2 = 6.93E-06   
+dw       = '1.15E-07+ddw_rnwaa'  
*+vc1     = 1.23E-02                vc2   = 8.92E-05  
+jc1a     = -2.80E-03              jc1b   = 2.66E-07    
+jc2a     = -3.10E-08              jc2b   = 3.21E-13
+rvc1     = 'jc1a+jc1b/l'          rvc2   =  '(jc2a+jc2b/l)/l' 
+weff     = 'w-2*dw'  
+tcoef(temper)     = '1.0+(temper-25.0)*(rtc1+rtc2*(temper-25.0))' 

D1    sub  n2 nwdioll area='weff*l/5' pj='weff+2*l/5'
R1    n2   na 'rsh*l/4/weff*tcoef(temper)*min(max(1.0+rvc1*v(n2,n1)+rvc2*v(n2,n1)*v(n2,n1), 0.85), 1.15)' 
D2    sub  na nwdioll area='weff*l/5' pj='2*l/5'
R2    na   nb 'rsh*l/4/weff*tcoef(temper)*min(max(1.0+rvc1*v(n2,n1)+rvc2*v(n2,n1)*v(n2,n1), 0.85), 1.15)' 
D3    sub  nb nwdioll area='weff*l/5' pj='2*l/5'
R3    nb   nc 'rsh*l/4/weff*tcoef(temper)*min(max(1.0+rvc1*v(n2,n1)+rvc2*v(n2,n1)*v(n2,n1), 0.85), 1.15)' 
D4    sub  nc nwdioll area='weff*l/5' pj='2*l/5'
R4    nc   n1 'rsh*l/4/weff*tcoef(temper)*min(max(1.0+rvc1*v(n2,n1)+rvc2*v(n2,n1)*v(n2,n1), 0.85), 1.15)' 
D5    sub  n1 nwdioll area='weff*l/5' pj='weff+2*l/5'  
.ends rnwaa_ckt  
************************************************************************************  
*        Silicide N+ diffusion resistor subcircuit netlist                         *  
************************************************************************************ 
.subckt rndif_ckt n2 n1 sub l=lr w=wr  
.param  
+rsh      = '14.131+drsh_rndif'    rtc1   = 2.00E-03       rtc2 = -3.43E-08   
+dw       = '-9.80E-09+ddw_rndif'  
*+vc1     = 6.53E-05               vc2   = 9.68E-05  
+jc1a     = 6.24E-05              jc1b   = 6.25E-10    
+jc2a     = 1.08E-08              jc2b   = 1.16E-12
+rvc1     = 'jc1a+jc1b/l'         rvc2   = '(jc2a+jc2b/l)/l' 
+weff     = 'w-2*dw' 
+tcoef(temper)     = '1.0+(temper-25.0)*(rtc1+rtc2*(temper-25.0))' 

D1    sub  n2 ndio12ll area='weff*l/5' pj='weff+2*l/5'
R1    n2   na 'rsh*l/4/weff*tcoef(temper)*min(1.0+rvc1*v(n2,n1)+rvc2*v(n2,n1)*v(n2,n1), 1.12)' 
D2    sub  na ndio12ll area='weff*l/5' pj='2*l/5'
R2    na   nb 'rsh*l/4/weff*tcoef(temper)*min(1.0+rvc1*v(n2,n1)+rvc2*v(n2,n1)*v(n2,n1), 1.12)' 
D3    sub  nb ndio12ll area='weff*l/5' pj='2*l/5'
R3    nb   nc 'rsh*l/4/weff*tcoef(temper)*min(1.0+rvc1*v(n2,n1)+rvc2*v(n2,n1)*v(n2,n1), 1.12)' 
D4    sub  nc ndio12ll area='weff*l/5' pj='2*l/5'
R4    nc   n1 'rsh*l/4/weff*tcoef(temper)*min(1.0+rvc1*v(n2,n1)+rvc2*v(n2,n1)*v(n2,n1), 1.12)' 
D5    sub  n1 ndio12ll area='weff*l/5' pj='weff+2*l/5'  
.ends rndif_ckt  
************************************************************************************  
*      Non-silicide N+ diffusion resistor subcircuit netlist                       *  
************************************************************************************ 
.subckt rndifsab_ckt n2 n1 sub l=lr w=wr  
.param  
+rsh      = '115.60+drsh_rndifsab'  rtc1   = 1.43E-03       rtc2 = 8.07E-07   
+dw       = '7.78E-09+ddw_rndifsab'   dl   = -1.88E-07
*+vc1     = 5.02E-04                 vc2   = 5.34E-03  
+jc1a     = 4.08E-04                jc1b   = 6.03E-10    
+jc2a     = 1.75E-08                jc2b   = 6.17E-14
+rvc1     = 'jc1a+jc1b/l'           rvc2   = '(jc2a+jc2b/l)/l' 
+weff     = 'w-2*dw'                leff   = 'l-2*dl'
+tcoef(temper)     = '1.0+(temper-25.0)*(rtc1+rtc2*(temper-25.0))' 

D1    sub  n2 ndio12ll area='weff*leff/5' pj='weff+2*leff/5'  
R1    n2   nb 'rsh*leff/4/weff*tcoef(temper)*min(1.0+rvc1*v(n2,n1)+rvc2*v(n2,n1)*v(n2,n1),1.12)'
D2    sub  nb ndio12ll area='weff*leff/5' pj='2*leff/5'
R2    nb   nc 'rsh*leff/4/weff*tcoef(temper)*min(1.0+rvc1*v(n2,n1)+rvc2*v(n2,n1)*v(n2,n1),1.12)'
D3    sub  nc ndio12ll area='weff*leff/5' pj='2*leff/5'
R3    nc   nd 'rsh*leff/4/weff*tcoef(temper)*min(1.0+rvc1*v(n2,n1)+rvc2*v(n2,n1)*v(n2,n1),1.12)'
D4    sub  nd ndio12ll area='weff*leff/5' pj='2*leff/5'
R4    nd   n1 'rsh*leff/4/weff*tcoef(temper)*min(1.0+rvc1*v(n2,n1)+rvc2*v(n2,n1)*v(n2,n1),1.12)'
D5    sub  n1 ndio12ll area='weff*leff/5' pj='weff+2*leff/5'  
.ends rndifsab_ckt   
************************************************************************************  
*        Silicide P+ diffusion resistor subcircuit netlist                         *  
************************************************************************************ 
.subckt rpdif_ckt n2 n1 sub l=lr w=wr  
.param  
+rsh      = '12.148+drsh_rpdif'      rtc1   = 2.49E-03       rtc2 = -7.68E-08   
+dw       = '-1.29E-08+ddw_rpdif'       
*+vc1     = -5.19E-06                vc2   = 2.39E-04  
+jc1a     = -7.61E-06               jc1b   = 4.49E-10    
+jc2a     = 2.59E-08                jc2b   = 1.35E-12
+rvc1     = 'jc1a+jc1b/l'           rvc2   = '(jc2a+jc2b/l)/l' 
+weff     = 'w-2*dw'   
+tcoef(temper)     = '1.0+(temper-25.0)*(rtc1+rtc2*(temper-25.0))' 

D1    n2  sub pdio12ll area='weff*l/5' pj='weff+2*l/5'
R1    n2   na 'rsh*l/4/weff*tcoef(temper)*min(1.0+rvc1*v(n2,n1)+rvc2*v(n2,n1)*v(n2,n1), 1.12)' 
D2    na  sub pdio12ll area='weff*l/5' pj='2*l/5'
R2    na   nb 'rsh*l/4/weff*tcoef(temper)*min(1.0+rvc1*v(n2,n1)+rvc2*v(n2,n1)*v(n2,n1), 1.12)' 
D3    nb  sub pdio12ll area='weff*l/5' pj='2*l/5'
R3    nb   nc 'rsh*l/4/weff*tcoef(temper)*min(1.0+rvc1*v(n2,n1)+rvc2*v(n2,n1)*v(n2,n1), 1.12)' 
D4    nc  sub pdio12ll area='weff*l/5' pj='2*l/5'
R4    nc   n1 'rsh*l/4/weff*tcoef(temper)*min(1.0+rvc1*v(n2,n1)+rvc2*v(n2,n1)*v(n2,n1), 1.12)' 
D5    n1  sub pdio12ll area='weff*l/5' pj='weff+2*l/5'   
.ends rpdif_ckt  
************************************************************************************  
*      Non-silicide P+ diffusion resistor subcircuit netlist                       *  
************************************************************************************ 
.subckt rpdifsab_ckt n2 n1 sub l=lr w=wr  
.param  
+rsh      = '259.00+drsh_rpdifsab'   rtc1   = 1.60E-03       rtc2 = 1.43E-06   
+dw       = '1.00E-09+ddw_rpdifsab'    dl   = -1.47E-07
*+vc1     = -5.08E-04                 vc2   = 2.97E-03  
+jc1a     = -8.98E-05                jc1b   = -2.70E-09    
+jc2a     = 1.45E-08                 jc2b   = 1.69E-14
+rvc1     = 'jc1a+jc1b/l'            rvc2   = '(jc2a+jc2b/l)/l' 
+weff     = 'w-2*dw'                 leff   = 'l-2*dl'
+tcoef(temper)     = '1.0+(temper-25.0)*(rtc1+rtc2*(temper-25.0))' 

D1    n2   sub pdio12ll area='weff*leff/5' pj='weff+2*leff/5'
R1    n2   na 'rsh*leff/4/weff*tcoef(temper)*min(1.0+rvc1*v(n2,n1)+rvc2*v(n2,n1)*v(n2,n1),1.11)'
D2    na   sub pdio12ll area='weff*leff/5' pj='2*leff/5'
R2    na   nb 'rsh*leff/4/weff*tcoef(temper)*min(1.0+rvc1*v(n2,n1)+rvc2*v(n2,n1)*v(n2,n1),1.11)'
D3    nb   sub pdio12ll area='weff*leff/5' pj='2*leff/5'
R3    nb   nc 'rsh*leff/4/weff*tcoef(temper)*min(1.0+rvc1*v(n2,n1)+rvc2*v(n2,n1)*v(n2,n1),1.11)'
D4    nc   sub pdio12ll area='weff*leff/5' pj='2*leff/5'
R4    nc   n1 'rsh*leff/4/weff*tcoef(temper)*min(1.0+rvc1*v(n2,n1)+rvc2*v(n2,n1)*v(n2,n1),1.11)'
D5    n1   sub pdio12ll area='weff*leff/5' pj='weff+2*leff/5'
.ends rpdifsab_ckt  
************************************************************************************  
*          Silicide N+ poly resistor subcircuit netlist                            *  
************************************************************************************ 
.subckt rnpo_ckt n2 n1 l=lr w=wr   
.param  
+rsh      = '13.405+drsh_rnpo'      rtc1   = 2.14E-03       rtc2 = -1.14E-07   
+dw       = '4.90E-09+ddw_rnpo'    
*+vc1     = 9.11E-05                vc2   = 5.16E-04  
+jc1a     = -7.37E-05              jc1b   = 3.60E-08    
+jc2a     = 3.75E-08               jc2b   = 8.48E-12
+rvc1     = 'jc1a+jc1b/l'          rvc2   = '(jc2a+jc2b/l)/l'          
+weff     = 'w-2*dw'
+tcoef(temper)     = '1.0+(temper-25.0)*(rtc1+rtc2*(temper-25.0))' 

R1 n2 n1 'rsh*l/weff*tcoef(temper)*min(1.0+rvc1*abs(v(n2,n1))+rvc2*v(n2,n1)*v(n2,n1), 1.26)'  
.ends rnpo_ckt  
************************************************************************************  
*          Silicide N+ poly resistor subcircuit netlist (three terminal)           *  
************************************************************************************ 
.subckt rnpo_3t_ckt n2 n1 sub l=lr w=wr   
.param  
+rsh      = '13.405+drsh_rnpo_3t'      rtc1   = 2.14E-03       rtc2 = -1.14E-07   
+dw       = '4.90E-09+ddw_rnpo_3t'    
*+vc1     = 9.11E-05                vc2   = 5.16E-04  
+jc1a     = -7.37E-05              jc1b   = 3.60E-08    
+jc2a     = 3.75E-08               jc2b   = 8.48E-12
+rvc1     = 'jc1a+jc1b/l'          rvc2   = '(jc2a+jc2b/l)/l'          
+weff     = 'w-2*dw'
+tcoef(temper)     = '1.0+(temper-25.0)*(rtc1+rtc2*(temper-25.0))' 
+cox      = 1.0117E-4             capsw   = 6.9120E-11

C1 n2 sub 'cox*weff*l/2+capsw*weff+capsw*l' 
R1 n2 n1 'rsh*l/weff*tcoef(temper)*min(1.0+rvc1*abs(v(n2,n1))+rvc2*v(n2,n1)*v(n2,n1), 1.26)'  
C2 n1 sub 'cox*weff*l/2+capsw*weff+capsw*l' 
.ends rnpo_3t_ckt  
************************************************************************************  
*        Non-silicide N+ poly resistor subcircuit netlist                          *  
************************************************************************************ 
.subckt rnposab_ckt n2 n1 l=lr w=wr  
.param  
+rsh      = '292.45+drsh_rnposab'   rtc1   = -2.49E-04           rtc2 = 4.67E-07   
+dw       = '2.27E-08+ddw_rnposab'    dl   = -1.29E-07
*+vc1     = -2.62E-05                vc2   = -4.98E-03  
+jc1a     = 1.94E-04                jc1b   = -1.34E-09    
+jc2a     = -4.32E-09               jc2b   = -8.87E-14
+rvc1     = 'jc1a+jc1b/l'           rvc2   = '(jc2a+jc2b/l)/l' 
+weff     = 'w-2*dw'                leff   = 'l-2*dl'
+tcoef(temper)     = '1.0+(temper-25.0)*(rtc1+rtc2*(temper-25.0))' 

R1    n2 n1 'rsh*leff/weff*tcoef(temper)*max(1.0+rvc1*abs(v(n2,n1))+rvc2*v(n2,n1)*v(n2,n1),0.834)'
.ends rnposab_ckt  
************************************************************************************  
*        Non-silicide N+ poly resistor subcircuit netlist (three terminal)         *  
************************************************************************************ 
.subckt rnposab_3t_ckt n2 n1 sub l=lr w=wr  
.param  
+rsh      = '292.45+drsh_rnposab_3t'   rtc1   = -2.49E-04           rtc2 = 4.67E-07   
+dw       = '2.27E-08+ddw_rnposab_3t'    dl   = -1.29E-07
*+vc1     = -2.62E-05                vc2   = -4.98E-03  
+jc1a     = 1.94E-04                jc1b   = -1.34E-09    
+jc2a     = -4.32E-09               jc2b   = -8.87E-14
+rvc1     = 'jc1a+jc1b/l'           rvc2   = '(jc2a+jc2b/l)/l' 
+weff     = 'w-2*dw'                leff   = 'l-2*dl'
+tcoef(temper)     = '1.0+(temper-25.0)*(rtc1+rtc2*(temper-25.0))' 
+cox      = 1.0117E-4              capsw   = 6.9120E-11

C1    n2 sub 'cox*weff*leff/2+capsw*weff+capsw*leff' 
R1    n2 n1 'rsh*leff/weff*tcoef(temper)*max(1.0+rvc1*abs(v(n2,n1))+rvc2*v(n2,n1)*v(n2,n1),0.834)'
C2    n1 sub 'cox*weff*leff/2+capsw*weff+capsw*leff'
.ends rnposab_3t_ckt  
************************************************************************************  
*          Silicide P+ poly resistor subcircuit netlist                            *  
************************************************************************************ 
.subckt rppo_ckt n2 n1 l=lr w=wr   
.param  
+rsh      = '12.420+drsh_rppo'      rtc1   = 2.47E-03       rtc2 = -9.28E-08   
+dw       = '4E-09+ddw_rppo'      
*+vc1     = 1.45E-04                vc2   = 6.53E-04  
+jc1a     = -1.02E-04              jc1b   = 5.40E-08    
+jc2a     = 4.89E-08               jc2b   = 1.06E-11
+rvc1     = 'jc1a+jc1b/l'          rvc2   = '(jc2a+jc2b/l)/l'          
+weff     = 'w-2*dw' 
+tcoef(temper)     = '1.0+(temper-25.0)*(rtc1+rtc2*(temper-25.0))' 

R1 n2 n1 'rsh*l/weff*tcoef(temper)*min(1.0+rvc1*abs(v(n2,n1))+rvc2*v(n2,n1)*v(n2,n1), 1.22)'  
.ends rppo_ckt  
************************************************************************************  
*          Silicide P+ poly resistor subcircuit netlist (three terminal)           *  
************************************************************************************ 
.subckt rppo_3t_ckt n2 n1 sub l=lr w=wr   
.param  
+rsh      = '12.420+drsh_rppo_3t'      rtc1   = 2.47E-03       rtc2 = -9.28E-08   
+dw       = '4E-09+ddw_rppo_3t'      
*+vc1     = 1.45E-04                vc2   = 6.53E-04  
+jc1a     = -1.02E-04              jc1b   = 5.40E-08    
+jc2a     = 4.89E-08               jc2b   = 1.06E-11
+rvc1     = 'jc1a+jc1b/l'          rvc2   = '(jc2a+jc2b/l)/l'          
+weff     = 'w-2*dw' 
+tcoef(temper)     = '1.0+(temper-25.0)*(rtc1+rtc2*(temper-25.0))' 
+cox      = 1.0117E-4              capsw   = 6.9120E-11

C1 n2 sub 'cox*weff*l/2+capsw*weff+capsw*l' 
R1 n2 n1 'rsh*l/weff*tcoef(temper)*min(1.0+rvc1*abs(v(n2,n1))+rvc2*v(n2,n1)*v(n2,n1), 1.22)'  
C2 n1 sub 'cox*weff*l/2+capsw*weff+capsw*l'
.ends rppo_3t_ckt 
************************************************************************************  
*        Non-silicide P+ poly resistor subcircuit netlist                          *  
************************************************************************************ 
.subckt rpposab_ckt n2 n1 l=lr w=wr  
.param  
+rsh      = '679.210+drsh_rpposab'   rtc1   = -3.04E-04       rtc2 = 5.33E-07   
+dw       = '2.79E-08+ddw_rpposab'    dl   = -1.00E-07
*+vc1     = -4.77E-04                vc2   = -1.69E-03  
+jc1a     = 1.29E-04                jc1b   = -3.91E-09    
+jc2a     = -3.37E-09               jc2b   = -2.73E-14
+rvc1     = 'jc1a+jc1b/l'           rvc2   = '(jc2a+jc2b/l)/l' 
+weff     = 'w-2*dw'                leff   = 'l-2*dl'
+tcoef(temper)     = '1.0+(temper-25.0)*(rtc1+rtc2*(temper-25.0))' 

R1    n2 n1 'rsh*leff/weff*tcoef(temper)*max(1.0+rvc1*abs(v(n2,n1))+rvc2*v(n2,n1)*v(n2,n1),0.892)'
.ends rpposab_ckt 
************************************************************************************  
*        Non-silicide P+ poly resistor subcircuit netlist (three terminal)         *  
************************************************************************************ 
.subckt rpposab_3t_ckt n2 n1 sub l=lr w=wr  
.param  
+rsh      = '679.210+drsh_rpposab_3t'   rtc1   = -3.04E-04       rtc2 = 5.33E-07   
+dw       = '2.79E-08+ddw_rpposab_3t'     dl   = -1.00E-07
*+vc1     = -4.77E-04                vc2   = -1.69E-03  
+jc1a     = 1.29E-04                jc1b   = -3.91E-09    
+jc2a     = -3.37E-09               jc2b   = -2.73E-14
+rvc1     = 'jc1a+jc1b/l'           rvc2   = '(jc2a+jc2b/l)/l' 
+weff     = 'w-2*dw'                leff   = 'l-2*dl'
+tcoef(temper)     = '1.0+(temper-25.0)*(rtc1+rtc2*(temper-25.0))' 
+cox      = 1.0117E-4              capsw   = 6.9120E-11

C1    n2 sub 'cox*weff*leff/2+capsw*weff+capsw*leff' 
R1    n2 n1 'rsh*leff/weff*tcoef(temper)*max(1.0+rvc1*abs(v(n2,n1))+rvc2*v(n2,n1)*v(n2,n1),0.892)'
C2    n1 sub 'cox*weff*leff/2+capsw*weff+capsw*leff'
.ends rpposab_3t_ckt 
*****************************************  
*          Metal 1 resistance           *  
*****************************************
.subckt rm1_ckt n2 n1 sub l=lr w=wr   
.param  
+rsh       = '0.1288+drsh_rm1'      rtc1  = 3.20E-03           rtc2  = 3.92E-07   
+dw        = '8.40E-09+ddw_rm1'     
*+vc1      = 0                       vc2  = 1.18E-03
+jc1a      = 0                      jc1b  = 0
+jc2a      = 1.69E-07               jc2b  = 1.38E-10
+rvc1      = 'jc1a+jc1b/l'          rvc2  = '(jc2a+jc2b/l)/l'          
+weff      = 'w-2*dw'              
+tcoef(temper)     = '1.0+(temper-25.0)*(rtc1+rtc2*(temper-25.0))' 
+cox       = 4.6333E-05            capsw  = 1.0044E-10


C1 n2 sub 'cox*weff*l/2+capsw*weff+capsw*l'    
R1 n2 n1 'rsh*l/weff*tcoef(temper)*min(1.0+rvc1*abs(v(n2,n1))+rvc2*v(n2,n1)*v(n2,n1), 1.1)'
C2 n1 sub 'cox*weff*l/2+capsw*weff+capsw*l'  
.ends rm1_ckt
*****************************************  
*          Metal 2 resistance           *  
*****************************************
.subckt rm2_ckt n2 n1 sub l=lr w=wr   
.param  
+rsh       = '0.0948+drsh_rm2'      rtc1  = 3.29E-03           rtc2  = 3.88E-07   
+dw        = '1.61E-08+ddw_rm2'     
*+vc1      = 0                       vc2  = 1.37E-03
+jc1a      = 0                      jc1b  = 0
+jc2a      = 2.85E-07               jc2b  = 1.64E-10
+rvc1      = 'jc1a+jc1b/l'          rvc2  = '(jc2a+jc2b/l)/l'          
+weff      = 'w-2*dw'              
+tcoef(temper)     = '1.0+(temper-25.0)*(rtc1+rtc2*(temper-25.0))' 
+cox       = 3.0000E-05            capsw  = 9.3210E-11

C1 n2 sub 'cox*weff*l/2+capsw*weff+capsw*l'    
R1 n2 n1 'rsh*l/weff*tcoef(temper)*min(1.0+rvc1*abs(v(n2,n1))+rvc2*v(n2,n1)*v(n2,n1), 1.1)'
C2 n1 sub 'cox*weff*l/2+capsw*weff+capsw*l'  
.ends rm2_ckt
*****************************************  
*          Metal 3 resistance           *  
*****************************************
.subckt rm3_ckt n2 n1 sub l=lr w=wr   
.param  
+rsh       = '0.0948+drsh_rm3'      rtc1  = 3.29E-03           rtc2  = 3.88E-07   
+dw        = '1.61E-08+ddw_rm3'     
*+vc1      = 0                       vc2  = 1.37E-03
+jc1a      = 0                      jc1b  = 0
+jc2a      = 2.85E-07               jc2b  = 1.64E-10
+rvc1      = 'jc1a+jc1b/l'          rvc2  = '(jc2a+jc2b/l)/l'          
+weff      = 'w-2*dw'              
+tcoef(temper)     = '1.0+(temper-25.0)*(rtc1+rtc2*(temper-25.0))' 
+cox       = 2.1200E-05            capsw  = 9.2990E-11

C1 n2 sub 'cox*weff*l/2+capsw*weff+capsw*l'    
R1 n2 n1 'rsh*l/weff*tcoef(temper)*min(1.0+rvc1*abs(v(n2,n1))+rvc2*v(n2,n1)*v(n2,n1), 1.1)'
C2 n1 sub 'cox*weff*l/2+capsw*weff+capsw*l'  
.ends rm3_ckt
*****************************************  
*          Metal 4 resistance           *  
*****************************************
.subckt rm4_ckt n2 n1 sub l=lr w=wr   
.param  
+rsh       = '0.0948+drsh_rm4'      rtc1  = 3.29E-03           rtc2  = 3.88E-07   
+dw        = '1.61E-08+ddw_rm4'     
*+vc1      = 0                       vc2  = 1.37E-03
+jc1a      = 0                      jc1b  = 0
+jc2a      = 2.85E-07               jc2b  = 1.64E-10
+rvc1      = 'jc1a+jc1b/l'          rvc2  = '(jc2a+jc2b/l)/l'          
+weff      = 'w-2*dw'              
+tcoef(temper)     = '1.0+(temper-25.0)*(rtc1+rtc2*(temper-25.0))' 
+cox       = 1.6400E-05            capsw  = 9.2810E-11

C1 n2 sub 'cox*weff*l/2+capsw*weff+capsw*l'    
R1 n2 n1 'rsh*l/weff*tcoef(temper)*min(1.0+rvc1*abs(v(n2,n1))+rvc2*v(n2,n1)*v(n2,n1), 1.1)'
C2 n1 sub 'cox*weff*l/2+capsw*weff+capsw*l'  
.ends rm4_ckt
*****************************************  
*          Metal 5 resistance           *  
*****************************************
.subckt rm5_ckt n2 n1 sub l=lr w=wr   
.param  
+rsh       = '0.0948+drsh_rm5'      rtc1  = 3.29E-03           rtc2  = 3.88E-07   
+dw        = '1.61E-08+ddw_rm5'     
*+vc1      = 0                       vc2  = 1.37E-03
+jc1a      = 0                      jc1b  = 0
+jc2a      = 2.85E-07               jc2b  = 1.64E-10
+rvc1      = 'jc1a+jc1b/l'          rvc2  = '(jc2a+jc2b/l)/l'          
+weff      = 'w-2*dw'              
+tcoef(temper)     = '1.0+(temper-25.0)*(rtc1+rtc2*(temper-25.0))' 
+cox       = 1.3300E-05            capsw  = 9.2730E-11

C1 n2 sub 'cox*weff*l/2+capsw*weff+capsw*l'    
R1 n2 n1 'rsh*l/weff*tcoef(temper)*min(1.0+rvc1*abs(v(n2,n1))+rvc2*v(n2,n1)*v(n2,n1), 1.1)'
C2 n1 sub 'cox*weff*l/2+capsw*weff+capsw*l'  
.ends rm5_ckt
*****************************************  
*          Metal 6 resistance           *  
*****************************************
.subckt rm6_ckt n2 n1 sub l=lr w=wr   
.param  
+rsh       = '0.0948+drsh_rm6'      rtc1  = 3.29E-03           rtc2  = 3.88E-07   
+dw        = '1.61E-08+ddw_rm6'     
*+vc1      = 0                       vc2  = 1.37E-03
+jc1a      = 0                      jc1b  = 0
+jc2a      = 2.85E-07               jc2b  = 1.64E-10
+rvc1      = 'jc1a+jc1b/l'          rvc2  = '(jc2a+jc2b/l)/l'          
+weff      = 'w-2*dw'              
+tcoef(temper)     = '1.0+(temper-25.0)*(rtc1+rtc2*(temper-25.0))' 
+cox       = 1.1300E-05            capsw  = 9.2740E-11

C1 n2 sub 'cox*weff*l/2+capsw*weff+capsw*l'    
R1 n2 n1 'rsh*l/weff*tcoef(temper)*min(1.0+rvc1*abs(v(n2,n1))+rvc2*v(n2,n1)*v(n2,n1), 1.1)'
C2 n1 sub 'cox*weff*l/2+capsw*weff+capsw*l'  
.ends rm6_ckt
*****************************************  
*          Metal 7 resistance           *  
*****************************************
.subckt rm7_ckt n2 n1 sub l=lr w=wr   
.param  
+rsh       = '0.0948+drsh_rm7'      rtc1  = 3.29E-03           rtc2  = 3.88E-07   
+dw        = '1.61E-08+ddw_rm7'     
*+vc1      = 0                       vc2  = 1.37E-03
+jc1a      = 0                      jc1b  = 0
+jc2a      = 2.85E-07               jc2b  = 1.64E-10
+rvc1      = 'jc1a+jc1b/l'          rvc2  = '(jc2a+jc2b/l)/l'          
+weff      = 'w-2*dw'              
+tcoef(temper)     = '1.0+(temper-25.0)*(rtc1+rtc2*(temper-25.0))' 
+cox       = 9.7400E-06            capsw  = 9.2710E-11

C1 n2 sub 'cox*weff*l/2+capsw*weff+capsw*l'    
R1 n2 n1 'rsh*l/weff*tcoef(temper)*min(1.0+rvc1*abs(v(n2,n1))+rvc2*v(n2,n1)*v(n2,n1), 1.1)'
C2 n1 sub 'cox*weff*l/2+capsw*weff+capsw*l'  
.ends rm7_ckt
*****************************************  
*          Metal 8 resistance           *  
*****************************************
.subckt rm8_ckt n2 n1 sub l=lr w=wr   
.param  
+rsh       = '0.0948+drsh_rm8'      rtc1  = 3.29E-03           rtc2  = 3.88E-07   
+dw        = '1.61E-08+ddw_rm8'     
*+vc1      = 0                       vc2  = 1.37E-03
+jc1a      = 0                      jc1b  = 0
+jc2a      = 2.85E-07               jc2b  = 1.64E-10
+rvc1      = 'jc1a+jc1b/l'          rvc2  = '(jc2a+jc2b/l)/l'          
+weff      = 'w-2*dw'              
+tcoef(temper)     = '1.0+(temper-25.0)*(rtc1+rtc2*(temper-25.0))' 
+cox       = 8.5800E-06            capsw  = 1.0211E-10

C1 n2 sub 'cox*weff*l/2+capsw*weff+capsw*l'    
R1 n2 n1 'rsh*l/weff*tcoef(temper)*min(1.0+rvc1*abs(v(n2,n1))+rvc2*v(n2,n1)*v(n2,n1), 1.1)'
C2 n1 sub 'cox*weff*l/2+capsw*weff+capsw*l'  
.ends rm8_ckt
*****************************************  
*        Top Metal 1 resistance         *  
*****************************************
.subckt rtm1_ckt n2 n1 sub l=lr w=wr   
.param  
+rsh       = '0.0180+drsh_rtm1'      rtc1  = 3.76E-03           rtc2  = 3.45E-07   
+dw        = '1.80E-08+ddw_rtm1'     
*+vc1      = 0                        vc2  = 7.98E-03
+jc1a      = 0                       jc1b  = 0
+jc2a      = 1.83E-06                jc2b  = 2.25E-10
+rvc1      = 'jc1a+jc1b/l'           rvc2  = '(jc2a+jc2b/l)/l'          
+weff      = 'w-2*dw'              
+tcoef(temper)     = '1.0+(temper-25.0)*(rtc1+rtc2*(temper-25.0))' 
+cox       = 6.8333E-06             capsw  = 1.1153E-10

C1 n2 sub 'cox*weff*l/2+capsw*weff+capsw*l'    
R1 n2 n1 'rsh*l/weff*tcoef(temper)*min(1.0+rvc1*abs(v(n2,n1))+rvc2*v(n2,n1)*v(n2,n1), 1.1)'
C2 n1 sub 'cox*weff*l/2+capsw*weff+capsw*l'  
.ends rtm1_ckt
*****************************************  
*        Top Metal 2 resistance         *  
*****************************************
.subckt rtm2_ckt n2 n1 sub l=lr w=wr   
.param  
+rsh       = '0.0180+drsh_rtm2'      rtc1  = 3.76E-03           rtc2  = 3.45E-07   
+dw        = '1.80E-08+ddw_rtm2'     
*+vc1      = 0                        vc2  = 7.98E-03
+jc1a      = 0                       jc1b  = 0
+jc2a      = 1.83E-06                jc2b  = 2.25E-10
+rvc1      = 'jc1a+jc1b/l'           rvc2  = '(jc2a+jc2b/l)/l'          
+weff      = 'w-2*dw'              
+tcoef(temper)     = '1.0+(temper-25.0)*(rtc1+rtc2*(temper-25.0))' 
+cox       = 5.2381E-06             capsw  = 1.1167E-10

C1 n2 sub 'cox*weff*l/2+capsw*weff+capsw*l'    
R1 n2 n1 'rsh*l/weff*tcoef(temper)*min(1.0+rvc1*abs(v(n2,n1))+rvc2*v(n2,n1)*v(n2,n1), 1.1)'
C2 n1 sub 'cox*weff*l/2+capsw*weff+capsw*l'  
.ends rtm2_ckt
*