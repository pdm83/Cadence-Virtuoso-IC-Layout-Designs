//* 
//* No part of this file can be released without the consent of SMIC.
//*
//*****************************************************************************************************************
//* SMIC 65nm Low Leakage 1P10M(1P9M, 1P8M, 1P7M, 1P6M) Salicide 1.2V/1.8V/2.5V SPICE model (for SPECTRE only) *
//*****************************************************************************************************************
//*
//* Release version    : 1.0
//*
//* Release date       : 09/30/2009
//*
//* Simulation tool    : Cadence spectre V6.2.1
//*
//*
//*  Resistor   :
//*        *------------------------------------------------* 
//*        |      Resistor      |  Resistor subckt          |
//*        *================================================*
//*        | N+ Diff SAB        |    rndifsab_ckt_rf        |
//*        *------------------------------------------------*
//*        | P+ Diff SAB        |    rpdifsab_ckt_rf        |
//*        *------------------------------------------------*
//*        | N+ poly SAB        |    rnposab_ckt_rf         |
//*        *------------------------------------------------*
//*        | p+ poly SAB        |    rpposab_ckt_rf         |
//*        *------------------------------------------------*
//*
simulator lang=spectre  insensitive=yes
ahdl_include "res_rf.va"

//************************************
//* Non-silicide N+ diffusion resistor
//************************************
//* l=length, w=width
subckt rndifsab_ckt_rf (port1 port2)
parameters l=0 w=0 devt=temp     
// +vc1 = 5.02E-04               vc2 = 5.34E-03
+ rjc1a = 4.08E-04             rjc1b = 6.03E-10
+ rjc2a = 1.75E-08             rjc2b = 6.17E-14
+  rtc1 = 1.43E-03              rtc2 = 8.07E-07
+    dw = 7.78E-09+ddw_rndifsab_rf   dl = -1.88E-07
+  tref = 25                     rsh = 115.60+drsh_rndifsab_rf

ls_rf    (1 port2) inductor    l=max((0.0050723*pwr(w*1e6,-1.1766)*pwr(l*1e6,-0.00054417*w*w*1e12+0.011442*w*1e6+2.9027))*1e-9, 1e-12)
cf_rf    (port1 1) capacitor   c=max((0.0135*w*1e6+0.173)*l*1e6*1e-15,1e-18)
rs_rf    (port1 1 port1 1) diffres_rf_hdl lr=l wr=w rtemp=devt etchl=dl etch=dw tc1=rtc1 tc2=rtc2 jc1a=rjc1a jc1b=rjc1b jc2a=rjc2a jc2b=rjc2b rsh0=rsh tnom=tref rmaxvcoef=1.12
rs2_rf   (1 port2) resistor    r=max(53.942*pwr(w*1e6,-1.6495)*exp((0.00093775*w*w*1e12-0.020084*w*1e6+0.29469)*l*1e6), 1e-3)
cf2_rf   (port1 4) capacitor   c=max(((0.0026416*pwr(w*1e6,1.9206))*l*1e6+(-0.045217*w*w*1e12-0.05115*w*1e6+0.53317))*1e-15,1e-18)
rs3_rf   (4 port2) resistor    r=max(220.86*pwr(l/w,1.6398),1e-3)
rsub1_rf (2 0)     resistor    r=max((29.664*w*1e6+19.21)*pwr(l*1e6,(0.0087308*w*w*1e12 - 0.18008*w*1e6 + 0.77314)), 1e-3)
csub1_rf (2 0)     capacitor   c=max((0.2353*l*1e6-0.8955)*1e-15,1e-18)
cox1_rf  (port1 2) capacitor   c=max(1.2814*pwr(l*w*1e12,0.85557)*1e-15, 1e-18)
rsub2_rf (3 0)     resistor    r=max((29.664*w*1e6+19.21)*pwr(l*1e6,(0.0087308*w*w*1e12 - 0.18008*w*1e6 + 0.77314)), 1e-3)
csub2_rf (3 0)     capacitor   c=max((0.2353*l*1e6-0.8955)*1e-15,1e-18)
cox2_rf  (port2 3) capacitor   c=max(1.2814*pwr(l*w*1e12,0.85557)*1e-15, 1e-18)
ends rndifsab_ckt_rf

//***********************************                                   
//*Non-silicide P+ Diffusion resistor               
//***********************************                      
//* l=length, w=width
subckt rpdifsab_ckt_rf (port1 port2)
parameters l=0 w=0 devt=temp   
// +vc1 = -5.08E-04               vc2 = 2.97E-03
+ rjc1a = -8.98E-05             rjc1b = -2.70E-09
+ rjc2a = 1.45E-08              rjc2b = 1.69E-14
+  rtc1 = 1.60E-03               rtc2 = 1.43E-06
+    dw = 1.00E-09+ddw_rpdifsab_rf    dl = -1.47E-07
+  tref = 25                      rsh = 259.00+drsh_rpdifsab_rf
 
ls_rf    (1 port2) inductor    l=max((0.0030891*pwr(w*1e6,-1.9837)+0.0000019)*pwr(l*1e6,3.2428)*1e-9, 1e-12)
cf_rf    (port1 1) capacitor   c=0.01*1e-15
rs_rf    (port1 1 port1 1) diffres_rf_hdl lr=l wr=w rtemp=devt etchl=dl etch=dw tc1=rtc1 tc2=rtc2 jc1a=rjc1a jc1b=rjc1b jc2a=rjc2a jc2b=rjc2b rsh0=rsh tnom=tref rmaxvcoef=1.11
rs2_rf   (1 port2) resistor    r=max(64.404*exp(0.174*l*1e6), 1e-3)
cf2_rf   (port1 4) capacitor   c=0.01*1e-15
rs3_rf   (4 port2) resistor    r=max(224.93*pwr(l/w,1.2419),1e-3)
rsub1_rf (2 0)     resistor    r=max(21.689*l/w+235.705, 1e-3)
csub1_rf (2 0)     capacitor   c=max((2.3549*w*1e6+6.2381)*1e-15,1e-18)
cox1_rf  (port1 2) capacitor   c=max(1.8043*pwr(l*w*1e12,0.587336)*1e-15, 1e-18)
rsub2_rf (3 0)     resistor    r=max(21.689*l/w+235.705, 1e-3)
csub2_rf (3 0)     capacitor   c=max((2.3549*w*1e6+6.2381)*1e-15,1e-18)
cox2_rf  (port2 3) capacitor   c=max(1.8043*pwr(l*w*1e12,0.587336)*1e-15, 1e-18)
ends rpdifsab_ckt_rf

//************************************             
//* Non-silicide N+ poly resistor             
//************************************             
//* l=length, w=width                          
subckt rnposab_ckt_rf (port1 port2)               
parameters l=0 w=0 devt=temp     
// +vc1 = -2.62E-05               vc2 = -4.98E-03
+ rjc1a = 1.94E-04              rjc1b = -1.34E-09
+ rjc2a = -4.32E-09             rjc2b = -8.87E-14
+  rtc1 = -2.49E-04              rtc2 = 4.67E-07
+    dw = 2.27E-08+ddw_rnposab_rf     dl = -1.29E-07
+  tref = 25                      rsh = 292.45+drsh_rnposab_rf

ls_rf    (1 port2) inductor    l=max(((0.0000071321*w*w*1e12-0.0001364*w*1e6+0.00075553)*pwr(l*1e6,0.0048517*w*w*1e12-0.067495*w*1e6+3.2819))*1e-9,1e-12)
cf_rf    (port1 1) capacitor   c=0.01*1e-15
rs_rf    (port1 1 port1 1) polyres_rf_hdl lr=l wr=w rtemp=devt etchl=dl etch=dw tc1=rtc1 tc2=rtc2 jc1a=rjc1a jc1b=rjc1b jc2a=rjc2a jc2b=rjc2b rsh0=rsh tnom=tref rminvcoef=0.834
rs2_rf   (1 port2) resistor    r=max(2619*exp(0.13262*l*1e6), 1e-3)
cf2_rf   (port1 4) capacitor   c=0.01*1e-15
rs3_rf   (4 port2) resistor    r=max(58.493*pwr(l/w,1.9161),1e-3)
rsub1_rf (2 0)     resistor    r=max(40.661*l/w+90.6515, 1e-3)
csub1_rf (2 0)     capacitor   c=max((0.012199*l*w*1e12+0.65835)*1e-15,1e-18)
cox1_rf  (port1 2) capacitor   c=max((0.063671*w*l*1e12 + 1.2)*1e-15, 1e-18)
rsub2_rf (3 0)     resistor    r=max(40.661*l/w+90.6515, 1e-3)
csub2_rf (3 0)     capacitor   c=max((0.012199*l*w*1e12+0.65835)*1e-15,1e-18)
cox2_rf  (port2 3) capacitor   c=max((0.063671*w*l*1e12 + 1.2)*1e-15, 1e-18)
ends rnposab_ckt_rf 
                                            
//************************************             
//* Non-silicide P+ poly resistor             
//************************************             
//* l=length, w=width                            
subckt rpposab_ckt_rf (port1 port2)               
parameters l=0 w=0 devt=temp      
// +vc1 = -4.77E-04               vc2 = -1.69E-03
+ rjc1a = 1.29E-04              rjc1b = -3.91E-09
+ rjc2a = -3.37E-09             rjc2b = -2.73E-14
+  rtc1 = -3.04E-04              rtc2 = 5.33E-07
+    dw = 2.79E-08+ddw_rpposab_rf     dl = -1.00E-07
+  tref = 25                      rsh = 679.210+drsh_rpposab_rf

ls_rf    (1 port2) inductor    l=max(((0.000044663*w*w*1e12-0.00090084*w*1e6+0.0057456)*pwr(l*1e6,0.00327*w*w*1e12-0.06319*w*1e6+3.2599))*1e-9, 1e-12)
cf_rf    (port1 1) capacitor   c=0.01*1e-15
rs_rf    (port1 1 port1 1) polyres_rf_hdl lr=l wr=w rtemp=devt etchl=dl etch=dw tc1=rtc1 tc2=rtc2 jc1a=rjc1a jc1b=rjc1b jc2a=rjc2a jc2b=rjc2b rsh0=rsh tnom=tref rminvcoef=0.892
rs2_rf   (1 port2) resistor    r=max(7561.1*exp(0.0908*l*1e6), 1e-3)
cf2_rf   (port1 4) capacitor   c=0.01*1e-15
rs3_rf   (4 port2) resistor    r=max(150.5*pwr(l/w,2.4743),1e-3)
rsub1_rf (2 0)     resistor    r=max(93.7805*l/w+187.84, 1e-3)
csub1_rf (2 0)     capacitor   c=max((0.013751*l*w*1e12+1.066455)*1e-15,1e-18)
cox1_rf  (port1 2) capacitor   c=max(0.18301*pwr(l*w*1e12,0.82036)*1e-15, 1e-18)
rsub2_rf (3 0)     resistor    r=max(93.7805*l/w+187.84, 1e-3)
csub2_rf (3 0)     capacitor   c=max((0.013751*l*w*1e12+1.066455)*1e-15,1e-18)
cox2_rf  (port2 3) capacitor   c=max(0.18301*pwr(l*w*1e12,0.82036)*1e-15, 1e-18)
ends rpposab_ckt_rf 
