* 
* No part of this file can be released without the consent of SMIC.
*
* Note: SMIC recommends that users set VNTOL=1E-9 at .option for more smooth convergence.
*************************************************************************************************************
* SMIC 65nm Low Leakage 1P10M(1P9M, 1P8M, 1P7M, 1P6M) Salicide 1.2V/1.8V/2.5V SPICE model (for HSPICE only) * 
*************************************************************************************************************
*
* Release version    : 1.0
*
* Release date       : 09/30/2009
*
* Simulation tool    : Synopsys Star-HSPICE version 2006.09-SP1
*
*  Resistor   :
*        *--------------------------------------------------* 
*        | Resistor           |    Resistor subckt          |
*        *==================================================*
*        | N+ Diff SAB        |    rndifsab_ckt_rf          | 
*        *--------------------------------------------------*
*        | P+ Diff SAB        |    rpdifsab_ckt_rf          |
*        *--------------------------------------------------*
*        | N+ poly SAB        |    rnposab_ckt_rf           |
*        *--------------------------------------------------*
*        | p+ poly SAB        |    rpposab_ckt_rf           |
*        *--------------------------------------------------*
*
**************************************                                   
* Non-silicide N+ Diffusion resistor *              
**************************************                      
.subckt rndifsab_ckt_rf port1 port2 l=l_rf w=w_rf 
.param
+rsh      = '115.60+drsh_rndifsab_rf'  rtc1   = 1.43E-03       rtc2 = 8.07E-07   
+dw       = '7.78E-09+ddw_rndifsab_rf'   dl   = -1.88E-07
*+vc1     = 5.02E-04                 vc2   = 5.34E-03  
+jc1a     = 4.08E-04                jc1b   = 6.03E-10    
+jc2a     = 1.75E-08                jc2b   = 6.17E-14
+rvc1     = 'jc1a+jc1b/l'           rvc2   = '(jc2a+jc2b/l)/l' 
+weff     = 'w-2*dw'                leff   = 'l-2*dl'
+tcoef(temper)     = '1.0+(temper-25.0)*(rtc1+rtc2*(temper-25.0))' 
Ls_rf 1 port2    'max((0.0050723*pwr(w*1e6,-1.1766)*pwr(l*1e6,-0.00054417*w*w*1e12+0.011442*w*1e6+2.9027))*1e-9, 1e-12)'
Cf_rf port1 1    'max((0.0135*w*1e6+0.173)*l*1e6*1e-15,1e-18)'
Rs_rf port1 1      'rsh*leff/weff*tcoef(temper)*min(1.0+rvc1*v(port1,1)+rvc2*v(port1,1)*v(port1,1),1.12)'
Rs2_rf 1 port2   'max(53.942*pwr(w*1e6,-1.6495)*exp((0.00093775*w*w*1e12-0.020084*w*1e6+0.29469)*l*1e6), 1e-3)'
Cf2_rf port1 4   'max(((0.0026416*pwr(w*1e6,1.9206))*l*1e6+(-0.045217*w*w*1e12-0.05115*w*1e6+0.53317))*1e-15,1e-18)'
Rs3_rf 4 port2   'max(220.86*pwr(l/w,1.6398),1e-3)'
Rsub1_rf 2 0     'max((29.664*w*1e6+19.21)*pwr(l*1e6,(0.0087308*w*w*1e12 - 0.18008*w*1e6 + 0.77314)), 1e-3)'
Csub1_rf 2 0     'max((0.2353*l*1e6-0.8955)*1e-15,1e-18)'
Cox1_rf port1 2  'max(1.2814*pwr(l*w*1e12,0.85557)*1e-15, 1e-18)' 
Rsub2_rf 3 0     'max((29.664*w*1e6+19.21)*pwr(l*1e6,(0.0087308*w*w*1e12 - 0.18008*w*1e6 + 0.77314)), 1e-3)'
Csub2_rf 3 0     'max((0.2353*l*1e6-0.8955)*1e-15,1e-18)'
Cox2_rf port2 3  'max(1.2814*pwr(l*w*1e12,0.85557)*1e-15, 1e-18)' 
.ends rndifsab_ckt_rf
**************************************                                   
* Non-silicide P+ Diffusion resistor *               
**************************************                      
.subckt rpdifsab_ckt_rf port1 port2 l=l_rf w=w_rf 
.param
+rsh      = '259.00+drsh_rpdifsab_rf'   rtc1   = 1.60E-03       rtc2 = 1.43E-06   
+dw       = '1.00E-09+ddw_rpdifsab_rf'    dl   = -1.47E-07
*+vc1     = -5.08E-04                 vc2   = 2.97E-03  
+jc1a     = -8.98E-05                jc1b   = -2.70E-09    
+jc2a     = 1.45E-08                 jc2b   = 1.69E-14
+rvc1     = 'jc1a+jc1b/l'            rvc2   = '(jc2a+jc2b/l)/l' 
+weff     = 'w-2*dw'                 leff   = 'l-2*dl'
+tcoef(temper)     = '1.0+(temper-25.0)*(rtc1+rtc2*(temper-25.0))' 
Ls_rf 1 port2    'max((0.0030891*pwr(w*1e6,-1.9837)+0.0000019)*pwr(l*1e6,3.2428)*1e-9, 1e-12)' 
Cf_rf port1 1    '0.01*1e-15'
Rs_rf port1 1      'rsh*leff/weff*tcoef(temper)*min(1.0+rvc1*v(port1,1)+rvc2*v(port1,1)*v(port1,1),1.11)'
Rs2_rf 1 port2   'max(64.404*exp(0.174*l*1e6), 1e-3)'
Cf2_rf port1 4   '0.01*1e-15'
Rs3_rf 4 port2   'max(224.93*pwr(l/w,1.2419),1e-3)'
Rsub1_rf 2 0     'max(21.689*l/w+235.705, 1e-3)'
Csub1_rf 2 0     'max((2.3549*w*1e6+6.2381)*1e-15,1e-18)'
Cox1_rf port1 2  'max(1.8043*pwr(l*w*1e12,0.587336)*1e-15, 1e-18)'
Rsub2_rf 3 0     'max(21.689*l/w+235.705, 1e-3)'
Csub2_rf 3 0     'max((2.3549*w*1e6+6.2381)*1e-15,1e-18)'
Cox2_rf port2 3  'max(1.8043*pwr(l*w*1e12,0.587336)*1e-15, 1e-18)'
.ends rpdifsab_ckt_rf
*********************************                                   
* Non-silicide N+ Poly resistor *               
*********************************                      
.subckt rnposab_ckt_rf port1 port2 l=l_rf w=w_rf 
.param
+rsh      = '292.45+drsh_rnposab_rf'   rtc1   = -2.49E-04           rtc2 = 4.67E-07   
+dw       = '2.27E-08+ddw_rnposab_rf'    dl   = -1.29E-07
*+vc1     = -2.62E-05                vc2   = -4.98E-03  
+jc1a     = 1.94E-04                jc1b   = -1.34E-09    
+jc2a     = -4.32E-09               jc2b   = -8.87E-14
+rvc1     = 'jc1a+jc1b/l'           rvc2   = '(jc2a+jc2b/l)/l' 
+weff     = 'w-2*dw'                leff   = 'l-2*dl'
+tcoef(temper)     = '1.0+(temper-25.0)*(rtc1+rtc2*(temper-25.0))'
Ls_rf 1 port2    'max(((0.0000071321*w*w*1e12-0.0001364*w*1e6+0.00075553)*pwr(l*1e6,0.0048517*w*w*1e12-0.067495*w*1e6+3.2819))*1e-9,1e-12)' 
Cf_rf port1 1    '0.01*1e-15'
Rs_rf port1 1    'rsh*leff/weff*tcoef(temper)*max(1.0+rvc1*abs(v(port1,1))+rvc2*v(port1,1)*v(port1,1),0.834)'
Rs2_rf 1 port2   'max(2619*exp(0.13262*l*1e6), 1e-3)'
Cf2_rf port1 4   '0.01*1e-15'
Rs3_rf 4 port2   'max(58.493*pwr(l/w,1.9161),1e-3)'
Rsub1_rf 2 0     'max(40.661*l/w+90.6515, 1e-3)'
Csub1_rf 2 0     'max((0.012199*l*w*1e12+0.65835)*1e-15,1e-18)'
Cox1_rf port1 2  'max((0.063671*w*l*1e12 + 1.2)*1e-15, 1e-18)'  
Rsub2_rf 3 0     'max(40.661*l/w+90.6515, 1e-3)'
Csub2_rf 3 0     'max((0.012199*l*w*1e12+0.65835)*1e-15,1e-18)'
Cox2_rf port2 3  'max((0.063671*w*l*1e12 + 1.2)*1e-15, 1e-18)' 
.ends rnposab_ckt_rf
*********************************                                   
* Non-silicide P+ Poly resistor *               
*********************************                      
.subckt rpposab_ckt_rf port1 port2 l=l_rf w=w_rf 
.param
+rsh      = '679.210+drsh_rpposab_rf'   rtc1   = -3.04E-04       rtc2 = 5.33E-07   
+dw       = '2.79E-08+ddw_rpposab_rf'    dl   = -1.00E-07
*+vc1     = -4.77E-04                vc2   = -1.69E-03  
+jc1a     = 1.29E-04                jc1b   = -3.91E-09    
+jc2a     = -3.37E-09               jc2b   = -2.73E-14
+rvc1     = 'jc1a+jc1b/l'           rvc2   = '(jc2a+jc2b/l)/l' 
+weff     = 'w-2*dw'                leff   = 'l-2*dl'
+tcoef(temper)     = '1.0+(temper-25.0)*(rtc1+rtc2*(temper-25.0))' 
Ls_rf 1 port2    'max(((0.000044663*w*w*1e12-0.00090084*w*1e6+0.0057456)*pwr(l*1e6,0.00327*w*w*1e12-0.06319*w*1e6+3.2599))*1e-9, 1e-12)' 
Cf_rf port1 1    '0.01*1e-15'
Rs_rf port1 1    'rsh*leff/weff*tcoef(temper)*max(1.0+rvc1*abs(v(port1,1))+rvc2*v(port1,1)*v(port1,1),0.892)'
Rs2_rf 1 port2   'max(7561.1*exp(0.0908*l*1e6), 1e-3)'
Cf2_rf port1 4   '0.01*1e-15'
Rs3_rf 4 port2   'max(150.5*pwr(l/w,2.4743),1e-3)'
Rsub1_rf 2 0     'max(93.7805*l/w+187.84, 1e-3)'
Csub1_rf 2 0     'max((0.013751*l*w*1e12+1.066455)*1e-15,1e-18)'
Cox1_rf port1 2  'max(0.18301*pwr(l*w*1e12,0.82036)*1e-15, 1e-18)'  
Rsub2_rf 3 0     'max(93.7805*l/w+187.84, 1e-3)'
Csub2_rf 3 0     'max((0.013751*l*w*1e12+1.066455)*1e-15,1e-18)'
Cox2_rf port2 3  'max(0.18301*pwr(l*w*1e12,0.82036)*1e-15, 1e-18)' 
.ends rpposab_ckt_rf
