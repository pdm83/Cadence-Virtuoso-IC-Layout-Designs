***hspice Model Format 
** library ind_diff 
** * 
** * no part of this file can be released without the consent of smic. 
** * 
** ****************************************************************************************** 
** *         smic 0.065um mixed signal 1p8m 1.2v*1.8*2.5v spice model (for hspice only)         * 
** ****************************************************************************************** 
** * 
** * release version    : 0.1 
** * 
** * release date       : Mar.*30*2009 
** * 
** * simulation tool    : Synopsys Star-HSPICE version 2008.09-SP1 
** * 
***  Inductor   : 
***    *--------------------------------------*--------------------*--------------------*---------------------* 
***    |  Turn & Radius  | Turn=3,rin=30~90um | Turn=4,rin=30~90um | Turn=5,rin=30~90um | Turn=6,rin=30~90um  | 
***    *--------------------------------------*--------------------*--------------------*---------------------* 
***    |                 |   ind_diff_t3r30   |   ind_diff_t4r30   |   ind_diff_t5r30   |   ind_diff_t6r30    | 
***    *                 ---------------------*--------------------*--------------------*---------------------* 
***    |                 |   ind_diff_t3r40   |   ind_diff_t4r40   |   ind_diff_t5r40   |   ind_diff_t6r40    | 
***    *                 ---------------------*--------------------*--------------------* --------------------*       
***    |                 |   ind_diff_t3r50   |   ind_diff_t4r50   |   ind_diff_t5r50   |   ind_diff_t6r50    | 
***    *   Model Name    ---------------------*--------------------*--------------------*---------------------* 
***    |                 |   ind_diff_t3r60   |   ind_diff_t4r60   |   ind_diff_t5r60   |   ind_diff_t6r60    | 
***    *                 ---------------------*--------------------*--------------------*---------------------* 
***    |                 |   ind_diff_t3r70   |   ind_diff_t4r70   |   ind_diff_t5r70   |   ind_diff_t6r70    | 
***    *                 ---------------------*--------------------*--------------------*---------------------* 
***    |                 |   ind_diff_t3r80   |   ind_diff_t4r80   |   ind_diff_t5r80   |   ind_diff_t6r80    | 
***    *                 ---------------------*--------------------*--------------------*---------------------* 
***    |                 |   ind_diff_t3r90   |   ind_diff_t4r90   |   ind_diff_t5r90   |   ind_diff_t6r90    | 
***    *--------------------------------------*--------------------*--------------------*---------------------* 
***   
***  
***     
*********************************************** 
*** 0.065um Three Port Differential Inductor 
*********************************************** 
.subckt ind_diff_t3r30 PLUS MINUS CT 
** *********************************************************************************** 
** *********************************************************************************** 
*****PLUS=port1(TM1**TM2), MINUS=port2(TM1**TM2), CT=Center Tap(M1**M2**M3)***** 
*****0.065um differential octagonal inductor two port equivalent circuit Single model***** 
*****n=3, w=8um, s=2.0um, TM1**TM2 inductor, rin=30um***** 
*****rin= inner radius; n= turns; w=width; s=spacing***** 
*****spacing is fixed at 2.0um, width is fixed at 8um and n is fixed at 3***** 
** *********************************************************************************** 
** *********************************************************************************** 
rs1 PLUS D 0.802 
ls1 D C 0.279e-9 
rsk1 PLUS D1 0.41 
lsk1 D1 D 0.060e-9 
ls2 C E 0.278e-9 
rs2 E MINUS 1.05 
rsk2 E E1 0.49 
lsk2 E1 MINUS 0.06e-9 
Kml1 ls1 ls2 0.585 
cs PLUS MINUS 13.57e-15 
lshort C F 0.226e-9 
rshort F CT 0.345 
rssk F F1 7.64 
lssk F1 CT 0.7565e-9 
cox1 PLUS A 15.85e-15 
csub1 A 0 1.343e-15 
rsub1 A 0 1558.0 
cox2 MINUS B 15.85e-15 
csub2 B 0 1.343e-15 
rsub2 B 0 1558.0 
.ends ind_diff_t3r30 

.subckt ind_diff_t3r40 PLUS MINUS CT 
** *********************************************************************************** 
** *********************************************************************************** 
*****PLUS=port1(TM1**TM2), MINUS=port2(TM1**TM2), CT=Center Tap(M1**M2**M3)***** 
*****0.065um differential octagonal inductor two port equivalent circuit Single model***** 
*****n=3, w=8um, s=2.0um, TM1**TM2 inductor, rin=40um***** 
*****rin= inner redius; n= turns; w=width; s=spacing***** 
*****spacing is fixed at 2.0um, width is fixed at 8um and n is fixed at 3***** 
** *********************************************************************************** 
** *********************************************************************************** 
rs1 PLUS D 0.817 
ls1 D C 0.38e-9 
rsk1 PLUS D1 0.7 
lsk1 D1 D 0.099e-9 
ls2 C E 0.385e-9 
rs2 E MINUS 0.901 
rsk2 E E1 0.92 
lsk2 E1 MINUS 0.143e-9 
Kml1 ls1 ls2 0.585 
cs PLUS MINUS 25.65e-15 
lshort C F 0.216e-9 
rshort F CT 0.331 
rssk F F1 7.64 
lssk F1 CT 0.7565e-9 
cox1 PLUS A 19.81e-15 
csub1 A 0 3.793e-15 
rsub1 A 0 1386.0 
cox2 MINUS B 19.81e-15 
csub2 B 0 3.793e-15 
rsub2 B 0 1386.0 
.ends ind_diff_t3r40 

.subckt ind_diff_t3r50 PLUS MINUS CT 
** *********************************************************************************** 
** *********************************************************************************** 
*****PLUS=port1(TM1**TM2), MINUS=port2(TM1**TM2), CT=Center Tap(M1**M2**M3)***** 
*****0.065um differential octagonal inductor two port equivalent circuit Single model***** 
*****n=3, w=8um, s=2.0um, TM1**TM2 inductor, rin=50um***** 
*****rin= inner redius; n= turns; w=width; s=spacing***** 
*****spacing is fixed at 2.0um, width is fixed at 8um and n is fixed at 3***** 
** *********************************************************************************** 
** *********************************************************************************** 
rs1 PLUS D 0.91 
ls1 D C 0.48e-9 
rsk1 PLUS D1 0.69 
lsk1 D1 D 0.101e-9 
ls2 C E 0.49e-9 
rs2 E MINUS 0.9 
rsk2 E E1 0.67 
lsk2 E1 MINUS 0.13e-9 
Kml1 ls1 ls2 0.585 
cs PLUS MINUS 38.22e-15 
lshort C F 0.218e-9 
rshort F CT 0.430 
rssk F F1 7.64 
lssk F1 CT 0.7565e-9 
cox1 PLUS A 18.92e-15 
csub1 A 0 9.019e-15 
rsub1 A 0 1172.0 
cox2 MINUS B 18.92e-15 
csub2 B 0 9.019e-15 
rsub2 B 0 1172.0 
.ends ind_diff_t3r50 

.subckt ind_diff_t3r60 PLUS MINUS CT 
** *********************************************************************************** 
** *********************************************************************************** 
*****PLUS=port1(TM1**TM2), MINUS=port2(TM1**TM2), CT=Center Tap(M1**M2**M3)***** 
*****0.065um differential octagonal inductor two port equivalent circuit Single model***** 
*****n=3, w=8um, s=2.0um, TM1**TM2 inductor, rin=60um***** 
*****rin= inner redius; n= turns; w=width; s=spacing***** 
*****spacing is fixed at 2.0um, width is fixed at 8um and n is fixed at 3***** 
** *********************************************************************************** 
** *********************************************************************************** 
rs1 PLUS D 1.2 
ls1 D C 0.59e-9 
rsk1 PLUS D1 1.06 
lsk1 D1 D 0.14e-9 
ls2 C E 0.60e-9 
rs2 E MINUS 1.2 
rsk2 E E1 1.2 
lsk2 E1 MINUS 0.18e-9 
Kml1 ls1 ls2 0.585 
cs PLUS MINUS 41.59e-15 
lshort C F 0.203e-9 
rshort F CT 0.370 
rssk F F1 7.64 
lssk F1 CT 0.7565e-9 
cox1 PLUS A 23.97e-15 
csub1 A 0 20.21e-15 
rsub1 A 0 986.0 
cox2 MINUS B 23.97e-15 
csub2 B 0 20.26e-15 
rsub2 B 0 986.0 
.ends ind_diff_t3r60 

.subckt ind_diff_t3r70 PLUS MINUS CT 
** *********************************************************************************** 
** *********************************************************************************** 
*****PLUS=port1(TM1**TM2), MINUS=port2(TM1**TM2), CT=Center Tap(M1**M2**M3)***** 
*****0.065um differential octagonal inductor two port equivalent circuit Single model***** 
*****n=3, w=8um, s=2.0um, TM1**TM2 inductor, rin=70um***** 
*****rin= inner redius; n= turns; w=width; s=spacing***** 
*****spacing is fixed at 2.0um, width is fixed at 8um and n is fixed at 3***** 
** *********************************************************************************** 
** *********************************************************************************** 
rs1 PLUS D 1.3 
ls1 D C 0.71e-9 
rsk1 PLUS D1 1.55 
lsk1 D1 D 0.176e-9 
ls2 C E 0.71e-9 
rs2 E MINUS 1.2 
rsk2 E E1 0.92 
lsk2 E1 MINUS 0.155e-9 
Kml1 ls1 ls2 0.585 
cs PLUS MINUS 49.11e-15 
lshort C F 0.203e-9 
rshort F CT 0.430 
rssk F F1 7.64 
lssk F1 CT 0.7565e-9 
cox1 PLUS A 18.0e-15 
csub1 A 0 11.83e-15 
rsub1 A 0 886.0 
cox2 MINUS B 18.0e-15 
csub2 B 0 11.83e-15 
rsub2 B 0 886.0 
.ends ind_diff_t3r70 

.subckt ind_diff_t3r80 PLUS MINUS CT 
** *********************************************************************************** 
** *********************************************************************************** 
*****PLUS=port1(TM1**TM2), MINUS=port2(TM1**TM2), CT=Center Tap(M1**M2**M3)***** 
*****0.065um differential octagonal inductor two port equivalent circuit Single model***** 
*****n=3, w=8um, s=2.0um, TM1**TM2 inductor, rin=80um***** 
*****rin= inner redius; n= turns; w=width; s=spacing***** 
*****spacing is fixed at 2.0um, width is fixed at 8um and n is fixed at 3***** 
** *********************************************************************************** 
** *********************************************************************************** 
rs1 PLUS D 1.4 
ls1 D C 0.82e-9 
rsk1 PLUS D1 1.57 
lsk1 D1 D 0.2e-9 
ls2 C E 0.83e-9 
rs2 E MINUS 1.27 
rsk2 E E1 1.2 
lsk2 E1 MINUS 0.2e-9 
Kml1 ls1 ls2 0.585 
cs PLUS MINUS 54.06e-15 
lshort C F 0.192e-9 
rshort F CT 0.430 
rssk F F1 7.64 
lssk F1 CT 0.7565e-9 
cox1 PLUS A 18.54e-15 
csub1 A 0 10.46e-15 
rsub1 A 0 858.0 
cox2 MINUS B 18.54e-15 
csub2 B 0 10.46e-15 
rsub2 B 0 858.0 
.ends ind_diff_t3r80 

.subckt ind_diff_t3r90 PLUS MINUS CT 
** *********************************************************************************** 
** *********************************************************************************** 
*****PLUS=port1(TM1**TM2), MINUS=port2(TM1**TM2), CT=Center Tap(M1**M2**M3)***** 
*****0.065um differential octagonal inductor two port equivalent circuit Single model***** 
*****n=3, w=8um, s=2.0um, TM1**TM2 inductor, rin=90um***** 
*****rin= inner redius; n= turns; w=width; s=spacing***** 
*****spacing is fixed at 2.0um, width is fixed at 8um and n is fixed at 3***** 
** *********************************************************************************** 
** *********************************************************************************** 
rs1 PLUS D 1.84 
ls1 D C 0.948e-9 
rsk1 PLUS D1 2.11 
lsk1 D1 D 0.29e-9 
ls2 C E 0.948e-9 
rs2 E MINUS 1.62 
rsk2 E E1 1.34 
lsk2 E1 MINUS 0.2e-9 
Kml1 ls1 ls2 0.585 
cs PLUS MINUS 59.61e-15 
lshort C F 0.182e-9 
rshort F CT 0.430 
rssk F F1 7.64 
lssk F1 CT 0.93e-9 
cox1 PLUS A 14.96e-15 
csub1 A 0 4.871e-15 
rsub1 A 0 700.0 
cox2 MINUS B 14.96e-15 
csub2 B 0 4.871e-15 
rsub2 B 0 700.0 
.ends ind_diff_t3r90 

.subckt ind_diff_t4r30 PLUS MINUS CT 
** *********************************************************************************** 
** *********************************************************************************** 
*****PLUS=port1(TM1**TM2), MINUS=port2(TM1**TM2), CT=Center Tap(M1**M2**M3)***** 
*****0.065um differential octagonal inductor two port equivalent circuit Single model***** 
*****n=4, w=8um, s=2.0um, TM1**TM2 inductor, rin=30um***** 
*****rin= inner redius; n= turns; w=width; s=spacing***** 
*****spacing is fixed at 2.0um, width is fixed at 8um and n is fixed at 4***** 
** *********************************************************************************** 
** *********************************************************************************** 
rs1 PLUS D 1.86 
ls1 D C 0.49e-9 
rsk1 PLUS D1 1.48 
lsk1 D1 D 0.176e-9 
ls2 C E 0.48e-9 
rs2 E MINUS 1.69 
rsk2 E E1 0.63 
lsk2 E1 MINUS 0.123e-9 
Kml1 ls1 ls2 0.603 
cs PLUS MINUS 46.34e-15 
lshort C F 0.254e-9 
rshort F CT 0.69 
rssk F F1 4.5 
lssk F1 CT 0.064e-9 
cox1 PLUS A 17.73e-15 
csub1 A 0 10.8e-15 
rsub1 A 0 1372.0 
cox2 MINUS B 17.73e-15 
csub2 B 0 10.8e-15 
rsub2 B 0 1372.0 
.ends ind_diff_t4r30 

.subckt ind_diff_t4r40 PLUS MINUS CT 
** *********************************************************************************** 
** *********************************************************************************** 
*****PLUS=port1(TM1**TM2), MINUS=port2(TM1**TM2), CT=Center Tap(M1**M2**M3)***** 
*****0.065um differential octagonal inductor two port equivalent circuit Single model***** 
*****n=4, w=8um, s=2.0um, TM1**TM2 inductor, rin=40um***** 
*****rin= inner redius; n= turns; w=width; s=spacing***** 
*****spacing is fixed at 2.0um, width is fixed at 8um and n is fixed at 4***** 
** *********************************************************************************** 
** *********************************************************************************** 
rs1 PLUS D 1.98 
ls1 D C 0.65e-9 
rsk1 PLUS D1 1.26 
lsk1 D1 D 0.176e-9 
ls2 C E 0.66e-9 
rs2 E MINUS 1.76 
rsk2 E E1 0.8 
lsk2 E1 MINUS 0.148e-9 
Kml1 ls1 ls2 0.603 
cs PLUS MINUS 55.35e-15 
lshort C F 0.239e-9 
rshort F CT 0.697 
rssk F F1 4.5 
lssk F1 CT 0.064e-9 
cox1 PLUS A 14.96e-15 
csub1 A 0 9.379e-15 
rsub1 A 0 1000 
cox2 MINUS B 14.96e-15 
csub2 B 0 9.379e-15 
rsub2 B 0 1000 
.ends ind_diff_t4r40 

.subckt ind_diff_t4r50 PLUS MINUS CT 
** *********************************************************************************** 
** *********************************************************************************** 
*****PLUS=port1(TM1**TM2), MINUS=port2(TM1**TM2), CT=Center Tap(M1**M2**M3)***** 
*****0.065um differential octagonal inductor two port equivalent circuit Single model***** 
*****n=4, w=8um, s=2.0um, TM1**TM2 inductor, rin=50um***** 
*****rin= inner redius; n= turns; w=width; s=spacing***** 
*****spacing is fixed at 2.0um, width is fixed at 8um and n is fixed at 4***** 
** *********************************************************************************** 
** *********************************************************************************** 
rs1 PLUS D 1.98 
ls1 D C 0.83e-9 
rsk1 PLUS D1 2.18 
lsk1 D1 D 0.282e-9 
ls2 C E 0.84e-9 
rs2 E MINUS 1.78 
rsk2 E E1 1.06 
lsk2 E1 MINUS 0.197e-9 
Kml1 ls1 ls2 0.603 
cs PLUS MINUS 63.07e-15 
lshort C F 0.233e-9 
rshort F CT 0.9272 
rssk F F1 4.5 
lssk F1 CT 0.064e-9 
cox1 PLUS A 16.94e-15 
csub1 A 0 12.56e-15 
rsub1 A 0 828.0 
cox2 MINUS B 16.94e-15 
csub2 B 0 12.56e-15 
rsub2 B 0 828.0 
.ends ind_diff_t4r50 

.subckt ind_diff_t4r60 PLUS MINUS CT 
** *********************************************************************************** 
** *********************************************************************************** 
*****PLUS=port1(TM1**TM2), MINUS=port2(TM1**TM2), CT=Center Tap(M1**M2**M3)***** 
*****0.065um differential octagonal inductor two port equivalent circuit Single model***** 
*****n=4, w=8um, s=2.0um, TM1**TM2 inductor, rin=60um***** 
*****rin= inner redius; n= turns; w=width; s=spacing***** 
*****spacing is fixed at 2.0um, width is fixed at 8um and n is fixed at 4***** 
** *********************************************************************************** 
** *********************************************************************************** 
rs1 PLUS D 2.46 
ls1 D C 1.01e-9 
rsk1 PLUS D1 1.83 
lsk1 D1 D 0.22e-9 
ls2 C E 1.01e-9 
rs2 E MINUS 2.04 
rsk2 E E1 1.06 
lsk2 E1 MINUS 0.197e-9 
Kml1 ls1 ls2 0.603 
cs PLUS MINUS 73.47e-15 
lshort C F 0.23e-9 
rshort F CT 1.00 
rssk F F1 4.5 
lssk F1 CT 0.064e-9 
cox1 PLUS A 12.88e-15 
csub1 A 0 4.136e-15 
rsub1 A 0 860.0 
cox2 MINUS B 12.88e-15 
csub2 B 0 4.136e-15 
rsub2 B 0 860.0 
.ends ind_diff_t4r60 

.subckt ind_diff_t4r70 PLUS MINUS CT 
** *********************************************************************************** 
** *********************************************************************************** 
*****PLUS=port1(TM1**TM2), MINUS=port2(TM1**TM2), CT=Center Tap(M1**M2**M3)***** 
*****0.065um differential octagonal inductor two port equivalent circuit Single model***** 
*****n=4, w=8um, s=2.0um, TM1**TM2 inductor, rin=70um***** 
*****rin= inner redius; n= turns; w=width; s=spacing***** 
*****spacing is fixed at 2.0um, width is fixed at 8um and n is fixed at 4***** 
** *********************************************************************************** 
** *********************************************************************************** 
rs1 PLUS D 2.36 
ls1 D C 1.2e-9 
rsk1 PLUS D1 1.83 
lsk1 D1 D 0.239e-9 
ls2 C E 1.2e-9 
rs2 E MINUS 2.32 
rsk2 E E1 1.34 
lsk2 E1 MINUS 0.218e-9 
Kml1 ls1 ls2 0.603 
cs PLUS MINUS 81.88e-15 
lshort C F 0.231e-9 
rshort F CT 1.14 
rssk F F1 4.5 
lssk F1 CT 0.064e-9 
cox1 PLUS A 15.5e-15 
csub1 A 0 6.586e-15 
rsub1 A 0 728 
cox2 MINUS B 15.5e-15 
csub2 B 0 6.586e-15 
rsub2 B 0 728 
.ends ind_diff_t4r70 

.subckt ind_diff_t4r80 PLUS MINUS CT 
** *********************************************************************************** 
** *********************************************************************************** 
*****PLUS=port1(TM1**TM2), MINUS=port2(TM1**TM2), CT=Center Tap(M1**M2**M3)***** 
*****0.065um differential octagonal inductor two port equivalent circuit Single model***** 
*****n=4, w=8um, s=2.0um, TM1**TM2 inductor, rin=80um***** 
*****rin= inner redius; n= turns; w=width; s=spacing***** 
*****spacing is fixed at 2.0um, width is fixed at 8um and n is fixed at 4***** 
** *********************************************************************************** 
** *********************************************************************************** 
rs1 PLUS D 2.28 
ls1 D C 1.38e-9 
rsk1 PLUS D1 1.54 
lsk1 D1 D 0.268e-9 
ls2 C E 1.39e-9 
rs2 E MINUS 2.01 
rsk2 E E1 1.43 
lsk2 E1 MINUS 0.3e-9 
Kml1 ls1 ls2 0.603 
cs PLUS MINUS 89.41e-15 
lshort C F 0.222e-9 
rshort F CT 1.28 
rssk F F1 3.29 
lssk F1 CT 0.07e-9 
cox1 PLUS A 18.92e-15 
csub1 A 0 5.9e-15 
rsub1 A 0 672 
cox2 MINUS B 18.92e-15 
csub2 B 0 5.9e-15 
rsub2 B 0 672 
.ends ind_diff_t4r80 

.subckt ind_diff_t4r90 PLUS MINUS CT 
** *********************************************************************************** 
** *********************************************************************************** 
*****PLUS=port1(TM1**TM2), MINUS=port2(TM1**TM2), CT=Center Tap(M1**M2**M3)***** 
*****0.065um differential octagonal inductor two port equivalent circuit Single model***** 
*****n=4, w=8um, s=2.0um, TM1**TM2 inductor, rin=90um***** 
*****rin= inner redius; n= turns; w=width; s=spacing***** 
*****spacing is fixed at 2.0um, width is fixed at 8um and n is fixed at 4***** 
** *********************************************************************************** 
** *********************************************************************************** 
rs1 PLUS D 2.18 
ls1 D C 1.59e-9 
rsk1 PLUS D1 1.47 
lsk1 D1 D 0.261e-9 
ls2 C E 1.59e-9 
rs2 E MINUS 2.18 
rsk2 E E1 1.15 
lsk2 E1 MINUS 0.26e-9 
Kml1 ls1 ls2 0.603 
cs PLUS MINUS 96.54e-15 
lshort C F 0.218e-9 
rshort F CT 1.34 
rssk F F1 4.5 
lssk F1 CT 0.064e-9 
cox1 PLUS A 21.89e-15 
csub1 A 0 5.9e-15 
rsub1 A 0 700 
cox2 MINUS B 21.89e-15 
csub2 B 0 5.9e-15 
rsub2 B 0 700 
.ends ind_diff_t4r90 

.subckt ind_diff_t5r30 PLUS MINUS CT 
** *********************************************************************************** 
** *********************************************************************************** 
*****PLUS=port1(TM1**TM2), MINUS=port2(TM1**TM2), CT=Center Tap(M1**M2**M3)***** 
*****0.065um differential octagonal inductor two port equivalent circuit Single model***** 
*****n=5, w=8um, s=2.0um, TM1**TM2 inductor, rin=30um***** 
*****rin= inner redius; n= turns; w=width; s=spacing***** 
*****spacing is fixed at 2.0um, width is fixed at 8um and n is fixed at 5***** 
** *********************************************************************************** 
** *********************************************************************************** 
rs1 PLUS D 2.1 
ls1 D C 0.668e-9 
rsk1 PLUS D1 1.2 
lsk1 D1 D 0.22e-9 
ls2 C E 0.668e-9 
rs2 E MINUS 2.0 
rsk2 E E1 0.92 
lsk2 E1 MINUS 0.22e-9 
Kml1 ls1 ls2 0.915 
cs PLUS MINUS 68.91e-15 
lshort C F 0.31e-9 
rshort F CT 0.359 
rssk F F1 6.06 
lssk F1 CT 0.21e-9 
cox1 PLUS A 16.34e-15 
csub1 A 0 3.793e-15 
rsub1 A 0 1386.0 
cox2 MINUS B 16.34e-15 
csub2 B 0 3.793e-15 
rsub2 B 0 1386.0 
.ends ind_diff_t5r30 

.subckt ind_diff_t5r40 PLUS MINUS CT 
** *********************************************************************************** 
** *********************************************************************************** 
*****PLUS=port1(TM1**TM2), MINUS=port2(TM1**TM2), CT=Center Tap(M1**M2**M3)***** 
*****0.065um differential octagonal inductor two port equivalent circuit Single model***** 
*****n=5, w=8um, s=2.0um, TM1**TM2 inductor, rin=40um***** 
*****rin= inner redius; n= turns; w=width; s=spacing***** 
*****spacing is fixed at 2.0um, width is fixed at 8um and n is fixed at 5***** 
** *********************************************************************************** 
** *********************************************************************************** 
rs1 PLUS D 2.31 
ls1 D C 0.88e-9 
rsk1 PLUS D1 2.25 
lsk1 D1 D 0.338e-9 
ls2 C E 0.88e-9 
rs2 E MINUS 2.12 
rsk2 E E1 1.22 
lsk2 E1 MINUS 0.28e-9 
Kml1 ls1 ls2 0.915 
cs PLUS MINUS 80.79e-15 
lshort C F 0.328e-9 
rshort F CT 0.38 
rssk F F1 6.2 
lssk F1 CT 0.35e-9 
cox1 PLUS A 14.96e-15 
csub1 A 0 2.764e-15 
rsub1 A 0 1128.0 
cox2 MINUS B 14.96e-15 
csub2 B 0 2.764e-15 
rsub2 B 0 1128.0 
.ends ind_diff_t5r40 

.subckt ind_diff_t5r50 PLUS MINUS CT 
** *********************************************************************************** 
** *********************************************************************************** 
*****PLUS=port1(TM1**TM2), MINUS=port2(TM1**TM2), CT=Center Tap(M1**M2**M3)***** 
*****0.065um differential octagonal inductor two port equivalent circuit Single model***** 
*****n=5, w=8um, s=2.0um, TM1**TM2 inductor, rin=50um***** 
*****rin= inner redius; n= turns; w=width; s=spacing***** 
*****spacing is fixed at 2.0um, width is fixed at 8um and n is fixed at 5***** 
** *********************************************************************************** 
** *********************************************************************************** 
rs1 PLUS D 2.49 
ls1 D C 1.09e-9 
rsk1 PLUS D1 2.26 
lsk1 D1 D 0.35e-9 
ls2 C E 1.09e-9 
rs2 E MINUS 2.32 
rsk2 E E1 1.12 
lsk2 E1 MINUS 0.268e-9 
Kml1 ls1 ls2 0.915 
cs PLUS MINUS 92.78e-15 
lshort C F 0.327e-9 
rshort F CT 0.373 
rssk F F1 6.2 
lssk F1 CT 0.093e-9 
cox1 PLUS A 16.0e-15 
csub1 A 0 3.6e-15 
rsub1 A 0 900.0 
cox2 MINUS B 16.0e-15 
csub2 B 0 3.6e-15 
rsub2 B 0 900.0 
.ends ind_diff_t5r50 

.subckt ind_diff_t5r60 PLUS MINUS CT 
** *********************************************************************************** 
** *********************************************************************************** 
*****PLUS=port1(TM1**TM2), MINUS=port2(TM1**TM2), CT=Center Tap(M1**M2**M3)***** 
*****0.065um differential octagonal inductor two port equivalent circuit Single model***** 
*****n=5, w=8um, s=2.0um, TM1**TM2 inductor, rin=60um***** 
*****rin= inner redius; n= turns; w=width; s=spacing***** 
*****spacing is fixed at 2.0um, width is fixed at 8um and n is fixed at 5***** 
** *********************************************************************************** 
** *********************************************************************************** 
rs1 PLUS D 2.34 
ls1 D C 1.32e-9 
rsk1 PLUS D1 1.9 
lsk1 D1 D 0.35e-9 
ls2 C E 1.32e-9 
rs2 E MINUS 2.43 
rsk2 E E1 1.55 
lsk2 E1 MINUS 0.35e-9 
Kml1 ls1 ls2 0.915 
cs PLUS MINUS 104.9e-15 
lshort C F 0.338e-9 
rshort F CT 0.37 
rssk F F1 6.2 
lssk F1 CT 0.7e-9 
cox1 PLUS A 18.3e-15 
csub1 A 0 4.25443e-15 
rsub1 A 0 835.8 
cox2 MINUS B 18.3e-15 
csub2 B 0 4.25443e-15 
rsub2 B 0 835.8 
.ends ind_diff_t5r60 

.subckt ind_diff_t5r70 PLUS MINUS CT 
** *********************************************************************************** 
** *********************************************************************************** 
*****PLUS=port1(TM1**TM2), MINUS=port2(TM1**TM2), CT=Center Tap(M1**M2**M3)***** 
*****0.065um differential octagonal inductor two port equivalent circuit Single model***** 
*****n=5, w=8um, s=2.0um, TM1**TM2 inductor, rin=70um***** 
*****rin= inner redius; n= turns; w=width; s=spacing***** 
*****spacing is fixed at 2.0um, width is fixed at 8um and n is fixed at 5***** 
** *********************************************************************************** 
** *********************************************************************************** 
rs1 PLUS D 2.6 
ls1 D C 1.55e-9 
rsk1 PLUS D1 1.45 
lsk1 D1 D 0.29e-9 
ls2 C E 1.56e-9 
rs2 E MINUS 2.6 
rsk2 E E1 1.41 
lsk2 E1 MINUS 0.35e-9 
Kml1 ls1 ls2 0.915 
cs PLUS MINUS 116.7e-15 
lshort C F 0.35e-9 
rshort F CT 0.394 
rssk F F1 6.83 
lssk F1 CT 0.7e-9 
cox1 PLUS A 19.81e-15 
csub1 A 0 4.25443e-15 
rsub1 A 0 835.819 
cox2 MINUS B 19.81e-15 
csub2 B 0 4.25443e-15 
rsub2 B 0 835.819 
.ends ind_diff_t5r70 

.subckt ind_diff_t5r80 PLUS MINUS CT 
** *********************************************************************************** 
** *********************************************************************************** 
*****PLUS=port1(TM1**TM2), MINUS=port2(TM1**TM2), CT=Center Tap(M1**M2**M3)***** 
*****0.065um differential octagonal inductor two port equivalent circuit Single model***** 
*****n=5, w=8um, s=2.0um, TM1**TM2 inductor, rin=80um***** 
*****rin= inner redius; n= turns; w=width; s=spacing***** 
*****spacing is fixed at 2.0um, width is fixed at 8um and n is fixed at 5***** 
** *********************************************************************************** 
** *********************************************************************************** 
rs1 PLUS D 2.38 
ls1 D C 1.8e-9 
rsk1 PLUS D1 2.2 
lsk1 D1 D 0.52e-9 
ls2 C E 1.8e-9 
rs2 E MINUS 2.38 
rsk2 E E1 2.11 
lsk2 E1 MINUS 0.53e-9 
Kml1 ls1 ls2 0.915 
cs PLUS MINUS 126.0e-15 
lshort C F 0.35e-9 
rshort F CT 0.33 
rssk F F1 6.83 
lssk F1 CT 0.7e-9 
cox1 PLUS A 24.66e-15 
csub1 A 0 5.46e-15 
rsub1 A 0 749.72 
cox2 MINUS B 24.66e-15 
csub2 B 0 5.46e-15 
rsub2 B 0 749.72 
.ends ind_diff_t5r80 

.subckt ind_diff_t5r90 PLUS MINUS CT 
** *********************************************************************************** 
** *********************************************************************************** 
*****PLUS=port1(TM1**TM2), MINUS=port2(TM1**TM2), CT=Center Tap(M1**M2**M3)***** 
*****0.065um differential octagonal inductor two port equivalent circuit Single model***** 
*****n=5, w=8um, s=2.0um, TM1**TM2 inductor, rin=90um***** 
*****rin= inner redius; n= turns; w=width; s=spacing***** 
*****spacing is fixed at 2.0um, width is fixed at 8um and n is fixed at 5***** 
** *********************************************************************************** 
** *********************************************************************************** 
rs1 PLUS D 3.1 
ls1 D C 2.02e-9 
rsk1 PLUS D1 2.32 
lsk1 D1 D 0.42e-9 
ls2 C E 2.02e-9 
rs2 E MINUS 3.1 
rsk2 E E1 2.22 
lsk2 E1 MINUS 0.42e-9 
Kml1 ls1 ls2 0.915 
cs PLUS MINUS 140.6e-15 
lshort C F 0.35e-9 
rshort F CT 0.49 
rssk F F1 6.06 
lssk F1 CT 0.77e-9 
cox1 PLUS A 21.89e-15 
csub1 A 0 12.19e-15 
rsub1 A 0 775.0 
cox2 MINUS B 21.89e-15 
csub2 B 0 6.057e-15 
rsub2 B 0 775.0 
.ends ind_diff_t5r90 

.subckt ind_diff_t6r30 PLUS MINUS CT 
** *********************************************************************************** 
** *********************************************************************************** 
*****0.065um differential octagonal inductor two port equivalent circuit Single model***** 
*****n=6, w=8um, s=2.0um, TM1**TM2 inductor, rin=30um***** 
*****PLUS=port1, MINUS=port2, CT=Center Tap***** 
*****rin= inner redius; n= turns; w=width; s=spacing; t=conductor thickness***** 
*****spacing is fixed at 2.0um, width is fixed at 10um and n is fixed at 6***** 
** *********************************************************************************** 
** *********************************************************************************** 
rs1 PLUS D 2.43 
ls1 D C 0.999e-9 
rsk1 PLUS D1 1.48 
lsk1 D1 D 0.35e-9 
ls2 C E 1.0e-9 
rs2 E MINUS 2.39 
rsk2 E E1 1.2 
lsk2 E1 MINUS 0.35e-9 
Kml1 ls1 ls2 0.915 
cs PLUS MINUS 93.76e-15 
lshort C F 0.358e-9 
rshort F CT 0.55 
rssk F F1 6.441 
lssk F1 CT 0.21e-9 
cox1 PLUS A 33.77e-15 
csub1 A 0 6.586e-15 
rsub1 A 0 1628.0 
cox2 MINUS B 33.77e-15 
csub2 B 0 6.586e-15 
rsub2 B 0 1625.0 
.ends ind_diff_t6r30 

.subckt ind_diff_t6r40 PLUS MINUS CT 
** *********************************************************************************** 
** *********************************************************************************** 
*****0.065um differential octagonal inductor two port equivalent circuit Single model***** 
*****n=6, w=8um, s=2.0um, TM1**TM2 inductor, rin=40um***** 
*****PLUS=port1, MINUS=port2, CT=Center Tap***** 
*****rin= inner redius; n= turns; w=width; s=spacing; t=conductor thickness***** 
*****spacing is fixed at 2.0um, width is fixed at 10um and n is fixed at 6***** 
** *********************************************************************************** 
** *********************************************************************************** 
rs1 PLUS D 2.55 
ls1 D C 1.29e-9 
rsk1 PLUS D1 2.01 
lsk1 D1 D 0.47e-9 
ls2 C E 1.29e-9 
rs2 E MINUS 2.55 
rsk2 E E1 1.28 
lsk2 E1 MINUS 0.4e-9 
Kml1 ls1 ls2 0.915 
cs PLUS MINUS 109.0e-15 
lshort C F 0.40e-9 
rshort F CT 0.60 
rssk F F1 9.6 
lssk F1 CT 0.74e-9 
cox1 PLUS A 24.36e-15 
csub1 A 0 8.007e-15 
rsub1 A 0 1314.0 
cox2 MINUS B 24.36e-15 
csub2 B 0 8.007e-15 
rsub2 B 0 1314.0 
.ends ind_diff_t6r40 

.subckt ind_diff_t6r50 PLUS MINUS CT 
** *********************************************************************************** 
** *********************************************************************************** 
*****0.065um differential octagonal inductor two port equivalent circuit Single model***** 
*****n=6, w=8um, s=2.0um, TM1**TM2 inductor, rin=50um***** 
*****PLUS=port1, MINUS=port2, CT=Center Tap***** 
*****rin= inner redius; n= turns; w=width; s=spacing; t=conductor thickness***** 
*****spacing is fixed at 2.0um, width is fixed at 10um and n is fixed at 6***** 
** *********************************************************************************** 
** *********************************************************************************** 
rs1 PLUS D 2.57 
ls1 D C 1.6e-9 
rsk1 PLUS D1 2.39 
lsk1 D1 D 0.56e-9 
ls2 C E 1.6e-9 
rs2 E MINUS 2.54 
rsk2 E E1 1.83 
lsk2 E1 MINUS 0.49e-9 
Kml1 ls1 ls2 0.915 
cs PLUS MINUS 123.8e-15 
lshort C F 0.4e-9 
rshort F CT 0.88 
rssk F F1 8.94 
lssk F1 CT 0.58e-9 
cox1 PLUS A 27.53e-15 
csub1 A 0 11.49e-15 
rsub1 A 0 1258.0 
cox2 MINUS B 27.53e-15 
csub2 B 0 11.49e-15 
rsub2 B 0 1258.0 
.ends ind_diff_t6r50 

.subckt ind_diff_t6r60 PLUS MINUS CT 
** *********************************************************************************** 
** *********************************************************************************** 
*****0.065um differential octagonal inductor two port equivalent circuit Single model***** 
*****n=6, w=8um, s=2.0um, TM1**TM2 inductor, rin=60um***** 
*****PLUS=port1, MINUS=port2, CT=Center Tap***** 
*****rin= inner redius; n= turns; w=width; s=spacing; t=conductor thickness***** 
*****spacing is fixed at 2.0um, width is fixed at 10um and n is fixed at 6***** 
** *********************************************************************************** 
** *********************************************************************************** 
rs1 PLUS D 2.96 
ls1 D C 1.9e-9 
rsk1 PLUS D1 2.39 
lsk1 D1 D 0.56e-9 
ls2 C E 1.9e-9 
rs2 E MINUS 2.96 
rsk2 E E1 2.39 
lsk2 E1 MINUS 0.56e-9 
Kml1 ls1 ls2 0.915 
cs PLUS MINUS 139.7e-15 
lshort C F 0.42e-9 
rshort F CT 0.87 
rssk F F1 9.44 
lssk F1 CT 0.92e-9 
cox1 PLUS A 23.97e-15 
csub1 A 0 13.59e-15 
rsub1 A 0 958.0 
cox2 MINUS B 23.97e-15 
csub2 B 0 13.59e-15 
rsub2 B 0 958.0 
.ends ind_diff_t6r60 

.subckt ind_diff_t6r70 PLUS MINUS CT 
** *********************************************************************************** 
** *********************************************************************************** 
*****0.065um differential octagonal inductor two port equivalent circuit Single model***** 
*****n=6, w=8um, s=2.0um, TM1**TM2 inductor, rin=70um***** 
*****PLUS=port1, MINUS=port2, CT=Center Tap***** 
*****rin= inner redius; n= turns; w=width; s=spacing; t=conductor thickness***** 
*****spacing is fixed at 2.0um, width is fixed at 10um and n is fixed at 6***** 
** *********************************************************************************** 
** *********************************************************************************** 
rs1 PLUS D 2.82 
ls1 D C 2.22e-9 
rsk1 PLUS D1 2.75 
lsk1 D1 D 0.63e-9 
ls2 C E 2.22e-9 
rs2 E MINUS 2.82 
rsk2 E E1 2.54 
lsk2 E1 MINUS 0.7e-9 
Kml1 ls1 ls2 0.915 
cs PLUS MINUS 153.8e-15 
lshort C F 0.43e-9 
rshort F CT 0.985 
rssk F F1 9.86 
lssk F1 CT 2.3e-9 
cox1 PLUS A 31.0e-15 
csub1 A 0 19.12e-15 
rsub1 A 0 929.0 
cox2 MINUS B 31.0e-15 
csub2 B 0 19.12e-15 
rsub2 B 0 929.0 
.ends ind_diff_t6r70 

.subckt ind_diff_t6r80 PLUS MINUS CT 
** *********************************************************************************** 
** *********************************************************************************** 
*****0.065um differential octagonal inductor two port equivalent circuit Single model***** 
*****n=6, w=8um, s=2.0um, TM1**TM2 inductor, rin=80um***** 
*****PLUS=port1, MINUS=port2, CT=Center Tap***** 
*****rin= inner redius; n= turns; w=width; s=spacing; t=conductor thickness***** 
*****spacing is fixed at 2.0um, width is fixed at 10um and n is fixed at 6***** 
** *********************************************************************************** 
** *********************************************************************************** 
rs1 PLUS D 2.82 
ls1 D C 2.55e-9 
rsk1 PLUS D1 4.23 
lsk1 D1 D 0.99e-9 
ls2 C E 2.55e-9 
rs2 E MINUS 2.82 
rsk2 E E1 2.61 
lsk2 E1 MINUS 0.77e-9 
Kml1 ls1 ls2 0.915 
cs PLUS MINUS 166.6e-15 
lshort C F 0.45e-9 
rshort F CT 1.07 
rssk F F1 9.932 
lssk F1 CT 0.812e-9 
cox1 PLUS A 33.77e-15 
csub1 A 0 19.12e-15 
rsub1 A 0 838.0 
cox2 MINUS B 33.77e-15 
csub2 B 0 19.12e-15 
rsub2 B 0 838.0 
.ends ind_diff_t6r80 

.subckt ind_diff_t6r90 PLUS MINUS CT 
** *********************************************************************************** 
** *********************************************************************************** 
*****0.065um differential octagonal inductor two port equivalent circuit Single model***** 
*****n=6, w=8um, s=2.0um, TM1**TM2 inductor, rin=90um***** 
*****PLUS=port1, MINUS=port2, CT=Center Tap***** 
*****rin= inner redius; n= turns; w=width; s=spacing; t=conductor thickness***** 
*****spacing is fixed at 2.0um, width is fixed at 10um and n is fixed at 6***** 
** *********************************************************************************** 
** *********************************************************************************** 
rs1 PLUS D 3.1 
ls1 D C 2.9e-9 
rsk1 PLUS D1 4.3 
lsk1 D1 D 0.99e-9 
ls2 C E 2.9e-9 
rs2 E MINUS 3.1 
rsk2 E E1 2.96 
lsk2 E1 MINUS 0.92e-9 
Kml1 ls1 ls2 0.901 
cs PLUS MINUS 181.7e-15 
lshort C F 0.458e-9 
rshort F CT 1.02 
rssk F F1 10.7 
lssk F1 CT 0.85e-9 
cox1 PLUS A 33.77e-15 
csub1 A 0 13.57e-15 
rsub1 A 0 711.0 
cox2 MINUS B 33.77e-15 
csub2 B 0 13.57e-15 
rsub2 B 0 711.0 
.ends ind_diff_t6r90 

** endlibrary ind_diff 
